module sevenSeg (a1, a2, b, x);

input [3:0] a1;
input [3:0] a2;
input b;
output reg [7:0] x;

always @ (*) begin
  if (b) begin
    case (a1)
      4'b0000: x = 8'b1100_0000; //0
      4'b0001: x = 8'b1111_1001; //1
      4'b0010: x = 8'b1010_0100; //2
      4'b0011: x = 8'b1011_0000; //3
      4'b0100: x = 8'b1001_1001; //4
      4'b0101: x = 8'b1001_0010; //5
      4'b0110: x = 8'b1000_0010; //6
      4'b0111: x = 8'b1111_1000; //7
      4'b1000: x = 8'b1000_0000; //8
      4'b1001: x = 8'b1001_1000; //9
      4'b1010: x = 8'b1111_1111; //A
      4'b1011: x = 8'b1000_0011; //b
      4'b1100: x = 8'b1100_0110; //C
      4'b1101: x = 8'b1010_0001; //d
      4'b1110: x = 8'b1000_0110; //E
      4'b1111: x = 8'b1000_1110; //F
      default: x = 8'b1111_1111;
    endcase
  end else begin
    case (a2)
      4'b0000: x = 8'b1100_0000; //0
      4'b0001: x = 8'b1111_1001; //1
      4'b0010: x = 8'b1010_0100; //2
      4'b0011: x = 8'b1011_0000; //3
      4'b0100: x = 8'b1001_1001; //4
      4'b0101: x = 8'b1001_0010; //5
      4'b0110: x = 8'b1000_0010; //6
      4'b0111: x = 8'b1111_1000; //7
      4'b1000: x = 8'b1000_0000; //8
      4'b1001: x = 8'b1001_1000; //9
      4'b1010: x = 8'b1000_1000; //A
      4'b1011: x = 8'b1000_0011; //b
      4'b1100: x = 8'b1100_0110; //C
      4'b1101: x = 8'b1010_0001; //d
      4'b1110: x = 8'b1000_0110; //E
      4'b1111: x = 8'b1000_1110; //F
      default: x = 8'b1111_1111;
    endcase
  end
end

endmodule