module stateProcessor ();
  
endmodule