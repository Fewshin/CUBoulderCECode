`ifdef sim
  parameter divider = 32'10;
`else 
  parameter divider = 32'd1500000;
`endif